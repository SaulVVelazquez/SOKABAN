333333333
302111113
312111113
312111113
312111113
312111413
312111113
333333333