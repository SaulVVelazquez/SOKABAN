3333333333
3021111113
3121111113
3121111113
3121141113
3121111113
3121111113
3333333333