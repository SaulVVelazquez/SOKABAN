3333333333
3011111113
3111111213
3114111113
3121141113
3111241113
3111111713
3333333333