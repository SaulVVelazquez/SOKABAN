3333333333
3011111113
3111111113
3111111113
3112141113
3111111713
3111111113
3333333333