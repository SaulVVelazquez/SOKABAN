33333333333333333333
31111111114111111113
31111111112111111113
31111111111111111113
31111111110111111113
31111111111111111113
31111111112111111113
31111111111111111113